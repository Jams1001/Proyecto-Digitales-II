module tester1 (
    output reg clk, reset,
    output reg [11:0] fifo_out,
    output reg [3:0] almost_full, empty,
    input wire [3:0] push, pop, push_estr, pop_estr
);

always #1 clk <= ~clk;


initial begin 
    empty = 4'b0000;
    reset = 1;
    almost_full = 0;
    fifo_out = 0;
    clk = 0;
end

initial begin
    $dumpfile("arbitro1.vcd");
    $dumpvars;
    repeat(2) @(posedge clk);
    reset = 0;
    fifo_out <= 12'b000010010110;
    repeat(4) @(posedge clk);       
    fifo_out <= 12'b100011110000;
    repeat(2) @(posedge clk);
    empty <= 4'b0100;
    @(posedge clk);                  
    fifo_out <= 12'b110110100000;
    @(posedge clk);
    fifo_out <= 12'b110100011110;
    @(posedge clk);
    empty <= 0;
    fifo_out <= 12'b111000101001;
    @(posedge clk);
    fifo_out <= 12'b111000101001;
    @(posedge clk);
    fifo_out <= 12'b111100101001;
    @(posedge clk);
    almost_full[2] <= 1;
    fifo_out <= 12'b111100101001;
    repeat(5) @(posedge clk);
    $finish;
end
    
endmodule